`timescale 1ns / 1ps

module grid_points
	#(parameter pd = 12, parameter p = 22)(
	input wire clk,
	input wire valid,
	input wire [7:0] p0_idx_i,
	input wire [6*3+6*p-1:0] cur_data_real_i, cur_data_imag_i,
	output wire [7:0] p0_idx_o,
	output wire enhance_o, eval_done_o,
	output reg [34-1:0] p0_d0_0, p0_d1_0, p0_d2_0,
	output reg [34-1:0] p1_d0_0, p1_d1_0, p1_d2_0,
	output reg [34-1:0] p2_d0_0, p2_d1_0, p2_d2_0,
	output reg [34-1:0] p3_d0_0, p3_d1_0, p3_d2_0
	//output reg eval_done
	);
	wire [7:0] p0_idx_best;
	
	reg eval_done = 1'b0;
	reg [7:0] p0_idx = 8'b0; // index of initial simplex based on grid of start values
	reg [7:0] p0_idx_next = 8'b0;
	
	initial begin
		p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
		p0_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
		p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0
		
		p1_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
		p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
		p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0
		
		p2_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
		p2_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
		p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

		p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
		p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
		p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
	end
	
	reg [7:0] p0_cnt = 8'b11111011; // total p0 cnt 11111011 (251)
	
	//assign eval_done = (grd_pnt_idx == 8'b11111101) ? 1'b1 : 1'b0;
	//assign eval_done = ((grd_pnt_idx == grd_pnt_idx_i_next) & (finished_loop)) ? 1'b1 : 1'b0; // done at the step after enhance
	/*
	always @(*) begin
		$display("p0_idx: %d", p0_idx);
		$display("p0_idx_best: %d", p0_idx_best);
		$display("loop_done: %d", loop_done);
	end
	*/
	///*
	/*
	reg finished_loop = 1'b0;
	always @(posedge clk) begin
		if (valid) begin
			grd_pnt_idx = grd_pnt_idx + 1;
		end
		// last iteration enhances best start
		if (grd_pnt_idx == p0_cnt) begin
			$display("grd_pnt_idx == p0_cnt");
			grd_pnt_idx = grd_pnt_idx_i;
			finished_loop = 1'b1;
		end 
		if (eval_done) begin
			grd_pnt_idx = 8'b00000000;
			finished_loop = 1'b0;
		end
	end
	*/
	/*
	reg sleep = 1'b1;
	always @(cur_data_real_i, cur_data_imag_i) begin
		sleep = 1'b0;
		if (eval_done_i) begin
			sleep = 1'b1;
		end
	end
	*/
	/*
	reg flag = 1'b0;
	always @(cur_data_real_i, cur_data_imag_i) begin
		if (not busy) begin
			flag <= 1'b1;
		end
	end
	*/
	
	assign enhance_o = ((p0_idx == p0_idx_best) & loop_done) ? 1'b1 : 1'b0;
	// always block to decide next grid point index (next state)
	reg loop_done = 1'b0;
	always @(valid, cur_data_real_i, cur_data_imag_i) begin
		if (valid) begin
			if ((p0_idx == p0_idx_best) & loop_done) begin
				p0_idx_next <= 8'b0;
			end else if (p0_idx == p0_cnt) begin
				loop_done <= 1'b1;
				p0_idx_next <= p0_idx_best;
			end else if (~loop_done) begin
				p0_idx_next <= p0_idx + 1;
			end else begin
				p0_idx_next <= p0_idx_next;
			end
		end else begin
			p0_idx_next <= p0_idx_next;
		end
		if ((p0_idx == 8'b0) & loop_done) begin
			loop_done <= 1'b0;
			eval_done <= 1'b1;
		end else if (eval_done) begin
			eval_done <= 1'b0;
		end else begin
			eval_done <= eval_done;
		end
		/*
		// triggered by sensitivity list (change in cur_data_real_i, cur_data_imag_i)
		if (eval_done) begin
			eval_done <= 1'b0;
		end else begin
			eval_done <= 1'b1;
		end
		*/
	end
	
	always @(posedge clk) begin
		p0_idx <= p0_idx_next;
	end
	
	assign enhance_o = loop_done;
	assign p0_idx_best = p0_idx_i;
	assign p0_idx_o = p0_idx;
	assign eval_done_o = eval_done;
	
	always @(p0_idx) begin
		case(p0_idx)
		/*
			[[50, 450, 50], [50, 450, 100], [50, 450, 150], [50, 450, 200], [50, 450, 250], [50, 450, 300], [50, 500, 50], [50, 500, 100], 
			[50, 500, 150], [50, 500, 200], [50, 500, 250], [50, 500, 300], [50, 550, 50], [50, 550, 100], [50, 550, 150], [50, 550, 200], 
			[50, 550, 250], [50, 550, 300], [50, 600, 50], [50, 600, 100], [50, 600, 150], [50, 600, 200], [50, 600, 250], [50, 600, 300], 
			[50, 650, 50], [50, 650, 100], [50, 650, 150], [50, 650, 200], [50, 650, 250], [50, 650, 300], [50, 700, 50], [50, 700, 100], 
			[50, 700, 150], [50, 700, 200], [50, 700, 250], [50, 700, 300], [50, 750, 50], [50, 750, 100], [50, 750, 150], [50, 750, 200], 
			[50, 750, 250], [50, 750, 300], [100, 450, 50], [100, 450, 100], [100, 450, 150], [100, 450, 200], [100, 450, 250], [100, 450, 300], 
			[100, 500, 50], [100, 500, 100], [100, 500, 150], [100, 500, 200], [100, 500, 250], [100, 500, 300], [100, 550, 50], [100, 550, 100], 
			[100, 550, 150], [100, 550, 200], [100, 550, 250], [100, 550, 300], [100, 600, 50], [100, 600, 100], [100, 600, 150], [100, 600, 200], 
			[100, 600, 250], [100, 600, 300], [100, 650, 50], [100, 650, 100], [100, 650, 150], [100, 650, 200], [100, 650, 250], [100, 650, 300], 
			[100, 700, 50], [100, 700, 100], [100, 700, 150], [100, 700, 200], [100, 700, 250], [100, 700, 300], [100, 750, 50], [100, 750, 100], 
			[100, 750, 150], [100, 750, 200], [100, 750, 250], [100, 750, 300], [150, 450, 50], [150, 450, 100], [150, 450, 150], [150, 450, 200], 
			[150, 450, 250], [150, 450, 300], [150, 500, 50], [150, 500, 100], [150, 500, 150], [150, 500, 200], [150, 500, 250], [150, 500, 300], 
			[150, 550, 50], [150, 550, 100], [150, 550, 150], [150, 550, 200], [150, 550, 250], [150, 550, 300], [150, 600, 50], [150, 600, 100], 
			[150, 600, 150], [150, 600, 200], [150, 600, 250], [150, 600, 300], [150, 650, 50], [150, 650, 100], [150, 650, 150], [150, 650, 200], 
			[150, 650, 250], [150, 650, 300], [150, 700, 50], [150, 700, 100], [150, 700, 150], [150, 700, 200], [150, 700, 250], [150, 700, 300], 
			[150, 750, 50], [150, 750, 100], [150, 750, 150], [150, 750, 200], [150, 750, 250], [150, 750, 300], [200, 450, 50], [200, 450, 100], 
			[200, 450, 150], [200, 450, 200], [200, 450, 250], [200, 450, 300], [200, 500, 50], [200, 500, 100], [200, 500, 150], [200, 500, 200], 
			[200, 500, 250], [200, 500, 300], [200, 550, 50], [200, 550, 100], [200, 550, 150], [200, 550, 200], [200, 550, 250], [200, 550, 300], 
			[200, 600, 50], [200, 600, 100], [200, 600, 150], [200, 600, 200], [200, 600, 250], [200, 600, 300], [200, 650, 50], [200, 650, 100], 
			[200, 650, 150], [200, 650, 200], [200, 650, 250], [200, 650, 300], [200, 700, 50], [200, 700, 100], [200, 700, 150], [200, 700, 200], 
			[200, 700, 250], [200, 700, 300], [200, 750, 50], [200, 750, 100], [200, 750, 150], [200, 750, 200], [200, 750, 250], [200, 750, 300], 
			[250, 450, 50], [250, 450, 100], [250, 450, 150], [250, 450, 200], [250, 450, 250], [250, 450, 300], [250, 500, 50], [250, 500, 100], 
			[250, 500, 150], [250, 500, 200], [250, 500, 250], [250, 500, 300], [250, 550, 50], [250, 550, 100], [250, 550, 150], [250, 550, 200], 
			[250, 550, 250], [250, 550, 300], [250, 600, 50], [250, 600, 100], [250, 600, 150], [250, 600, 200], [250, 600, 250], [250, 600, 300], 
			[250, 650, 50], [250, 650, 100], [250, 650, 150], [250, 650, 200], [250, 650, 250], [250, 650, 300], [250, 700, 50], [250, 700, 100], 
			[250, 700, 150], [250, 700, 200], [250, 700, 250], [250, 700, 300], [250, 750, 50], [250, 750, 100], [250, 750, 150], [250, 750, 200], 
			[250, 750, 250], [250, 750, 300], [300, 450, 50], [300, 450, 100], [300, 450, 150], [300, 450, 200], [300, 450, 250], [300, 450, 300], 
			[300, 500, 50], [300, 500, 100], [300, 500, 150], [300, 500, 200], [300, 500, 250], [300, 500, 300], [300, 550, 50], [300, 550, 100], 
			[300, 550, 150], [300, 550, 200], [300, 550, 250], [300, 550, 300], [300, 600, 50], [300, 600, 100], [300, 600, 150], [300, 600, 200], 
			[300, 600, 250], [300, 600, 300], [300, 650, 50], [300, 650, 100], [300, 650, 150], [300, 650, 200], [300, 650, 250], [300, 650, 300], 
			[300, 700, 50], [300, 700, 100], [300, 700, 150], [300, 700, 200], [300, 700, 250], [300, 700, 300], [300, 750, 50], [300, 750, 100], 
			[300, 750, 150], [300, 750, 200], [300, 750, 250], [300, 750, 300]]
		*/
			// Initial point idx 0
			8'b00000000 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0
				
				p1_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0
				
				p2_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p2_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 1
			8'b00000001 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 2
			8'b00000010 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 3
			8'b00000011 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 4
			8'b00000100 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 5
			8'b00000101 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 6
			8'b00000110 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 7
			8'b00000111 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 8
			8'b00001000 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 9
			8'b00001001 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 10
			8'b00001010 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 11
			8'b00001011 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 12
			8'b00001100 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 13
			8'b00001101 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 14
			8'b00001110 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 15
			8'b00001111 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 16
			8'b00010000 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 17
			8'b00010001 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 18
			8'b00010010 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 19
			8'b00010011 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 20
			8'b00010100 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 21
			8'b00010101 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 22
			8'b00010110 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 23
			8'b00010111 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 24
			8'b00011000 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 25
			8'b00011001 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 26
			8'b00011010 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 27
			8'b00011011 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 28
			8'b00011100 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 29
			8'b00011101 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 30
			8'b00011110 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 31
			8'b00011111 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 32
			8'b00100000 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 33
			8'b00100001 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 34
			8'b00100010 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 35
			8'b00100011 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 36
			8'b00100100 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 37
			8'b00100101 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 38
			8'b00100110 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 39
			8'b00100111 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 40
			8'b00101000 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 41
			8'b00101001 : begin
				p0_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000000101000_0000000000000000000000; // 40.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000000110010_0000000000000000000000; // 50.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 42
			8'b00101010 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 43
			8'b00101011 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 44
			8'b00101100 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 45
			8'b00101101 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 46
			8'b00101110 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 47
			8'b00101111 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 48
			8'b00110000 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 49
			8'b00110001 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 50
			8'b00110010 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 51
			8'b00110011 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 52
			8'b00110100 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 53
			8'b00110101 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 54
			8'b00110110 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 55
			8'b00110111 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 56
			8'b00111000 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 57
			8'b00111001 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 58
			8'b00111010 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 59
			8'b00111011 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 60
			8'b00111100 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 61
			8'b00111101 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 62
			8'b00111110 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 63
			8'b00111111 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 64
			8'b01000000 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 65
			8'b01000001 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 66
			8'b01000010 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 67
			8'b01000011 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 68
			8'b01000100 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 69
			8'b01000101 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 70
			8'b01000110 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 71
			8'b01000111 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 72
			8'b01001000 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 73
			8'b01001001 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 74
			8'b01001010 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 75
			8'b01001011 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 76
			8'b01001100 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 77
			8'b01001101 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 78
			8'b01001110 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 79
			8'b01001111 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 80
			8'b01010000 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 81
			8'b01010001 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 82
			8'b01010010 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 83
			8'b01010011 : begin
				p0_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001010000_0000000000000000000000; // 80.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000001100100_0000000000000000000000; // 100.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 84
			8'b01010100 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 85
			8'b01010101 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 86
			8'b01010110 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 87
			8'b01010111 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 88
			8'b01011000 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 89
			8'b01011001 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 90
			8'b01011010 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 91
			8'b01011011 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 92
			8'b01011100 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 93
			8'b01011101 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 94
			8'b01011110 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 95
			8'b01011111 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 96
			8'b01100000 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 97
			8'b01100001 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 98
			8'b01100010 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 99
			8'b01100011 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 100
			8'b01100100 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 101
			8'b01100101 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 102
			8'b01100110 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 103
			8'b01100111 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 104
			8'b01101000 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 105
			8'b01101001 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 106
			8'b01101010 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 107
			8'b01101011 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 108
			8'b01101100 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 109
			8'b01101101 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 110
			8'b01101110 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 111
			8'b01101111 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 112
			8'b01110000 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 113
			8'b01110001 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 114
			8'b01110010 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 115
			8'b01110011 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 116
			8'b01110100 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 117
			8'b01110101 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 118
			8'b01110110 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 119
			8'b01110111 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 120
			8'b01111000 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 121
			8'b01111001 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 122
			8'b01111010 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 123
			8'b01111011 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 124
			8'b01111100 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 125
			8'b01111101 : begin
				p0_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000001111000_0000000000000000000000; // 120.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000010010110_0000000000000000000000; // 150.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 126
			8'b01111110 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 127
			8'b01111111 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 128
			8'b10000000 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 129
			8'b10000001 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 130
			8'b10000010 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 131
			8'b10000011 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 132
			8'b10000100 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 133
			8'b10000101 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 134
			8'b10000110 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 135
			8'b10000111 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 136
			8'b10001000 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 137
			8'b10001001 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 138
			8'b10001010 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 139
			8'b10001011 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 140
			8'b10001100 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 141
			8'b10001101 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 142
			8'b10001110 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 143
			8'b10001111 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 144
			8'b10010000 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 145
			8'b10010001 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 146
			8'b10010010 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 147
			8'b10010011 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 148
			8'b10010100 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 149
			8'b10010101 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 150
			8'b10010110 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 151
			8'b10010111 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 152
			8'b10011000 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 153
			8'b10011001 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 154
			8'b10011010 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 155
			8'b10011011 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 156
			8'b10011100 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 157
			8'b10011101 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 158
			8'b10011110 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 159
			8'b10011111 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 160
			8'b10100000 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 161
			8'b10100001 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 162
			8'b10100010 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 163
			8'b10100011 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 164
			8'b10100100 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 165
			8'b10100101 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 166
			8'b10100110 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 167
			8'b10100111 : begin
				p0_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000010100000_0000000000000000000000; // 160.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 168
			8'b10101000 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 169
			8'b10101001 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 170
			8'b10101010 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 171
			8'b10101011 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 172
			8'b10101100 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 173
			8'b10101101 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 174
			8'b10101110 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 175
			8'b10101111 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 176
			8'b10110000 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 177
			8'b10110001 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 178
			8'b10110010 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 179
			8'b10110011 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 180
			8'b10110100 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 181
			8'b10110101 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 182
			8'b10110110 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 183
			8'b10110111 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 184
			8'b10111000 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 185
			8'b10111001 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 186
			8'b10111010 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 187
			8'b10111011 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 188
			8'b10111100 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 189
			8'b10111101 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 190
			8'b10111110 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 191
			8'b10111111 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 192
			8'b11000000 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 193
			8'b11000001 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 194
			8'b11000010 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 195
			8'b11000011 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 196
			8'b11000100 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 197
			8'b11000101 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 198
			8'b11000110 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 199
			8'b11000111 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 200
			8'b11001000 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 201
			8'b11001001 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 202
			8'b11001010 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 203
			8'b11001011 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 204
			8'b11001100 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 205
			8'b11001101 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 206
			8'b11001110 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 207
			8'b11001111 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 208
			8'b11010000 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 209
			8'b11010001 : begin
				p0_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011001000_0000000000000000000000; // 200.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000011111010_0000000000000000000000; // 250.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 210
			8'b11010010 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 211
			8'b11010011 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 212
			8'b11010100 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 213
			8'b11010101 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 214
			8'b11010110 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 215
			8'b11010111 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000101101000_0000000000000000000000; // 360.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b000111000010_0000000000000000000000; // 450.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 216
			8'b11011000 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 217
			8'b11011001 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 218
			8'b11011010 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 219
			8'b11011011 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 220
			8'b11011100 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 221
			8'b11011101 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000110010000_0000000000000000000000; // 400.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b000111110100_0000000000000000000000; // 500.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 222
			8'b11011110 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 223
			8'b11011111 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 224
			8'b11100000 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 225
			8'b11100001 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 226
			8'b11100010 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 227
			8'b11100011 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000110111000_0000000000000000000000; // 440.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001000100110_0000000000000000000000; // 550.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 228
			8'b11100100 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 229
			8'b11100101 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 230
			8'b11100110 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 231
			8'b11100111 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 232
			8'b11101000 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 233
			8'b11101001 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b000111100000_0000000000000000000000; // 480.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 234
			8'b11101010 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 235
			8'b11101011 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 236
			8'b11101100 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 237
			8'b11101101 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 238
			8'b11101110 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 239
			8'b11101111 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001000001000_0000000000000000000000; // 520.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001010001010_0000000000000000000000; // 650.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 240
			8'b11110000 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 241
			8'b11110001 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 242
			8'b11110010 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 243
			8'b11110011 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 244
			8'b11110100 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 245
			8'b11110101 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001000110000_0000000000000000000000; // 560.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001010111100_0000000000000000000000; // 700.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			// Initial point idx 246
			8'b11110110 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000000110010_0000000000000000000000; // 50.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000000101000_0000000000000000000000; // 40.0
			end
			// Initial point idx 247
			8'b11110111 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000001100100_0000000000000000000000; // 100.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000001010000_0000000000000000000000; // 80.0
			end
			// Initial point idx 248
			8'b11111000 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000010010110_0000000000000000000000; // 150.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000001111000_0000000000000000000000; // 120.0
			end
			// Initial point idx 249
			8'b11111001 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000010100000_0000000000000000000000; // 160.0
			end
			// Initial point idx 250
			8'b11111010 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000011111010_0000000000000000000000; // 250.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000011001000_0000000000000000000000; // 200.0
			end
			// Initial point idx 251
			8'b11111011 : begin
				p0_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p0_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p0_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p1_d0_0 = 34'b000011110000_0000000000000000000000; // 240.0
				p1_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p1_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p2_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p2_d1_0 = 34'b001001011000_0000000000000000000000; // 600.0
				p2_d2_0 = 34'b000100101100_0000000000000000000000; // 300.0

				p3_d0_0 = 34'b000100101100_0000000000000000000000; // 300.0
				p3_d1_0 = 34'b001011101110_0000000000000000000000; // 750.0
				p3_d2_0 = 34'b000011110000_0000000000000000000000; // 240.0
			end
			default : begin
				p0_d0_0 = p0_d0_0;
				p0_d1_0 = p0_d1_0;
				p0_d2_0 = p0_d2_0;
				
				p1_d0_0 = p1_d0_0;
				p1_d1_0 = p1_d1_0;
				p1_d2_0 = p1_d2_0;
				
				p2_d0_0 = p2_d0_0;
				p2_d1_0 = p2_d1_0;
				p2_d2_0 = p2_d2_0;

				p3_d0_0 = p3_d0_0;
				p3_d1_0 = p3_d1_0; 
				p3_d2_0 = p3_d2_0;
			end
		endcase
	end
	
endmodule